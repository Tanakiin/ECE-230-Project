ieee
print("Hello VHDL");
