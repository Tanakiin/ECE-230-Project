ieee
print("Hello world")
