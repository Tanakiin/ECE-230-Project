-- main fucntion goes in HERE! ALU to be designed
